module clk_gen(
    input  wire   in_clk,
    input  wire   rst_n,
    output reg    c0,
    output reg    locked 
);
    
endmodule