module ex (
    input
);
    
endmodule