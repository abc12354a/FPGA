module spi(
    input  wire       clk,
    input  wire       rst_n,
    input  wire[15:0] data,
    input  wire       MISO,
    output wire       sck,
    output wire       cs_n,
    output wire       MOSI
);
    
endmodule